library verilog;
use verilog.vl_types.all;
entity Fibonacci_TB is
end Fibonacci_TB;
